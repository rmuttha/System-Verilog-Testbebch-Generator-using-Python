��m o d u l e   c o u n t e r   (  
         i n p u t   w i r e   c l k ,  
         i n p u t   w i r e   r e s _ n ,  
         o u t p u t   r e g   [ 7 : 0 ]   c n t _ o u t  
 ) ;  
  
         / /   I n t e r n a l   s i g n a l   f o r   c o u n t i n g  
         r e g   [ 7 : 0 ]   c o u n t ;  
  
         / /   S y n c h r o n o u s   c o u n t e r  
         a l w a y s   @ ( p o s e d g e   c l k   o r   n e g e d g e   r e s _ n )   b e g i n  
                 i f   ( ! r e s _ n )   b e g i n  
                         / /   R e s e t   c o n d i t i o n  
                         c o u n t   < =   8 ' b 0 ;  
                 e n d   e l s e   b e g i n  
                         / /   C o u n t   u p   c o n d i t i o n  
                         c o u n t   < =   c o u n t   +   1 ;  
                 e n d  
         e n d  
  
         / /   A s s i g n   o u t p u t  
         a s s i g n   c n t _ o u t   =   c o u n t ;  
  
 e n d m o d u l e  
 